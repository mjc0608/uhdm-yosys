package p;

typedef struct packed {
	integer r;
	integer th;
} C;

typedef struct packed {
	logic [63:0] [3:0] a;
} S;

endpackage

module top(input [3:0] x, output reg [3:0] y, z);

	integer k = '{0:1, default: 0};
	integer i = '{31:1, 23:1, 15:1, 8:1, default: 0};
	integer j = '{default: 1, 31:0};

	p::C l = '{th:170, r:1};

	logic [96:0] A = '{1, 2, 3};

	p::S m = '{64'h9, 64'h12, 64'h21};


	always_comb begin
		assert(32'b00000000000000000000000000000001 == k);
		assert(32'b10000000100000001000000100000000 == i);
		assert(32'b01111111111111111111111111111111 == j);

		assert(l == 64'b0000000000000000000000000000000100000000000000000000000010101010);
		assert(m == 192'b000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000100001);

		assert(A == 96'b000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000011);
	end

endmodule
